----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:39:53 04/01/2014 
-- Design Name: 
-- Module Name:    Ca2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Ca2 is
    Port ( valeur : in  STD_LOGIC_VECTOR (13 downto 0);
           sortie : out  STD_LOGIC_VECTOR (13 downto 0));
end Ca2;

architecture Behavioral of Ca2 is
signal temp : STD_LOGIC_VECTOR (13 downto 0);

begin
process(valeur)
begin
	temp <= not valeur + "00000000000001";
end process;
sortie <=temp;
end Behavioral;

